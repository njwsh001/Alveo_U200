`define BAR_ADDR_WIDTH      22
`define BAR_DATA_WIDTH      32
`define USER_ADDR_WIDTH     14
`define USER_DATA_WIDTH     32
`define REG_BLOCK_NUM       64


//below define module id
`define PCIE_WRAP_ID        0